module bus_intf(
);

endmodule